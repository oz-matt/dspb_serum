
module dspb_serum_qsys (
	clk_clk,
	reset_reset_n,
	pio_0_external_connection_export);	

	input		clk_clk;
	input		reset_reset_n;
	input	[7:0]	pio_0_external_connection_export;
endmodule
